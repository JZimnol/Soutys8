------------------------------------------------------------------------------------------------------------------------
--
-- Title   : Control unit
-- Design  : Soutys8
-- Author  : J.Zimnol
-- Company : AGH Krakow
--
------------------------------------------------------------------------------------------------------------------------
--
-- Description:
--     Control unit of the processor. Controls write_enable signals and MUX outputs.
--
------------------------------------------------------------------------------------------------------------------------

library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.softprocessor_constants.all;

--------------------------------------------------------------------------------
-- ENTITY CONTROL_UNIT
--------------------------------------------------------------------------------
entity Control_unit is
    port(
        in_SREG_flags       : in  std_logic_vector(7 downto 0);
        in_instruction_type : in  std_logic_vector(5 downto 0);

        out_control         : out std_logic_vector(CONTROL_BUS_WIDTH-1 downto 0)
    );
end Control_unit;

--------------------------------------------------------------------------------
-- ARCHITECTURE OF CONTROL_UNIT
--------------------------------------------------------------------------------
architecture Control_unit of Control_unit is
    signal s_control          : std_logic_vector(CONTROL_BUS_WIDTH-1 downto 0) := (others => '0');
    signal s_previous_alu_op  : std_logic_vector(4 downto 0) := (others => '0');

begin

    process (in_SREG_flags, in_instruction_type) begin
        case in_instruction_type is
            when INSTR_TYPE_ADD  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_ADD;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_AND  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_AND;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_ANDI =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_AND;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_BRCC =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= not in_SREG_flags(ALU_FLAG_C);
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_BRCS =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                --s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= in_SREG_flags(ALU_FLAG_C);
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_BREQ =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= in_SREG_flags(ALU_FLAG_Z);
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_BRNE =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= not in_SREG_flags(ALU_FLAG_Z);
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CBI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_MEMORY;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_MMIO;
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CBI;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '1';
            when INSTR_TYPE_CLC  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_C;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLH  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_H;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_I;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLN  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_N;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLS  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_S;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLT  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_T;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLV  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_V;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CLZ  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_CLEAR_Z;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_COM  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_NEG;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CP   =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SUB;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_CPI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SUB;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_DEC  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_DEC;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_EOR  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_XOR;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_IN   =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_MMIO;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_MEMORY;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_INC  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_INC;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_JMP  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_JUMP;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_LDI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_IMMEDIATE;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_LDS_MMIO  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_MMIO;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_MEMORY;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_LDS_SRAM  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_SRAM;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_MEMORY;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_LSL  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_LSL;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_LSR  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_LSR;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_MOV  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_REGISTER;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_NOP  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_OR   =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_OR;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_ORI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_OR;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_OUT  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_REGISTER;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '1';
            when INSTR_TYPE_POP  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_SRAM;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_MEMORY;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '1';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_PUSH =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_REGISTER;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '1';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_RJMP =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SBI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_MEMORY;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_MMIO;
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SBI;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '1';
            when INSTR_TYPE_SBR  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_OR;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEC  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_C;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEH  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_H;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEI  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_I;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEN  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_N;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SES  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_S;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SET  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_T;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEV  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_V;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SEZ  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SET_Z;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_STS_MMIO  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_MMIO;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_REGISTER;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_STS_SRAM  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_BRANCH;
                s_control(CONTROL_MUX_READ_DATA) <= MUX_READ_DATA_SRAM;
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_REGISTER;
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '1';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SUB  =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_REGISTER;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SUB;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when INSTR_TYPE_SUBI =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '1';
                s_control(CONTROL_MUX_SRC1_SEL) <= MUX_ALU_SRC1_SEL_REGISTER;
                s_control(CONTROL_MUX_SRC2_SEL) <= MUX_ALU_SRC2_SEL_IMMEDIATE;
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <= MUX_WRITE_DATA_SEL_ALU;
                s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <= ALU_OP_SUB;
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '1';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
            when others =>
                s_control(CONTROL_REGISTER_FILE_WRITE_ENABLE) <= '0';
                --s_control(CONTROL_MUX_SRC1_SEL) <=
                --s_control(CONTROL_MUX_SRC2_SEL) <=
                s_control(CONTROL_MUX_PC_SEL) <= MUX_PC_SEL_NEXT_INSTR;
                s_control(CONTROL_MUX_BRANCH_SEL) <= MUX_BRANCH_SEL_NO_BRANCH;
                --s_control(CONTROL_MUX_READ_DATA) <=
                --s_control(CONTROL_MUX_WRITE_DATA_UPPER downto CONTROL_MUX_WRITE_DATA_LOWER) <=
                --s_control(CONTROL_ALU_OP_TYPE_UPPER downto CONTROL_ALU_OP_TYPE_LOWER) <=
                s_control(CONTROL_ALU_MODIFY_FLAG_ENABLE) <= '0';
                s_control(CONTROL_SRAM_WRITE_ENABLE) <= '0';
                s_control(CONTROL_SRAM_PUSH_ENABLE)  <= '0';
                s_control(CONTROL_SRAM_POP_ENABLE)   <= '0';
                s_control(CONTROL_GPIO_WRITE_ENABLE) <= '0';
        end case;
    end process;

    out_control <= s_control;

end Control_unit;
